`include "sample_seq_item.sv"
`include "sample_seq_lib.sv"
`include "sample_driver.sv"
`include "sample_monitor.sv"
`include "sample_sequencer.sv"
`include "sample_agent.sv"
`include "sample_env.sv"
