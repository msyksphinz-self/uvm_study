class sample_sequencer extends uvm_sequencer #(sample_seq_item);
  `uvm_component_utils(sample_sequencer);
  `uvm_new_func
endclass // sample_sequencer
