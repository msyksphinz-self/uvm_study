`include "switch_item.sv"
`include "driver.sv"
`include "monitor.sv"
`include "sequence.sv"
`include "scoreboard.sv"
`include "agent.sv"
`include "env.sv"
