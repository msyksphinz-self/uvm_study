interface sample_if (input logic clk, rstz);
  logic [ 7: 0] addr, data;
  logic         valid;
endinterface // sample_if
