`include "arbiter2_rr_seq_item.sv"
`include "arbiter2_rr_driver.sv"
`include "arbiter2_rr_monitor.sv"
`include "arbiter2_rr_sequence.sv"
`include "arbiter2_rr_scoreboard.sv"
`include "arbiter2_rr_agent.sv"
`include "arbiter2_rr_env.sv"
